`timescale 1ns/1ps
`default_nettype none


module tb_control();

reg sysclk;
reg clk; 
reg clken;
reg clken_oop;
reg clear;
integer count;
localparam CLKLEN = 4;

always #1 sysclk <= ~sysclk ;

always @(posedge sysclk)
begin
  if (count == CLKLEN-1) 
  begin
     clk <= ~clk;
     if (clk == 0)
       clken <= 1;
     else
       clken_oop <= 1;
     count <= 0;
  end else begin
     count <= count + 1;
     clken <= 0;
     clken_oop <= 0;
  end
end  



reg [3:0] ir_opc;
wire [11:0] cword;
wire halt;

wire [3:0] CU_counter = CU.T;
wire [11:0] cword = CU.cword;

wire pc_en;
wire pc_incr;
wire mar_load;

wire ir_en, ir_load;
wire mem_en;
wire a_en;
wire a_load;

controlunit CU(
  .sysclk(sysclk),
  //.clken(clken),
  .clken_oop(clken_oop),
  .clear(clear),
  .ir_opc(ir_opc),
  .cword(cword),
  .halt(halt)
);

wire [5:0] T = CU.T;

initial begin
   clear = 1;
   sysclk = 0;
   count = 0;
   clk = 0;
   #1;
   clear = 0;
   #1;
   ir_opc = 4'b0000;
   
   #200;
   $finish;  
end

endmodule
